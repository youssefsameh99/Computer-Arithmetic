module sixty_four_bit_brentkung_direct(
    input  [63:0] A, B,
    input cin,
    output [63:0] sum,
    output cout
);

wire [63:0] g, p;
assign g = A & B;
assign p = A ^ B;

wire [64:0] C;
assign C[0] = cin;

wire G0_0, P0_0;
wire G0_1, P0_1;
wire G0_2, P0_2;
wire G0_3, P0_3;
wire G0_4, P0_4;
wire G0_5, P0_5;
wire G0_6, P0_6;
wire G0_7, P0_7;
wire G0_8, P0_8;
wire G0_9, P0_9;
wire G0_10, P0_10;
wire G0_11, P0_11;
wire G0_12, P0_12;
wire G0_13, P0_13;
wire G0_14, P0_14;
wire G0_15, P0_15;
wire G0_16, P0_16;
wire G0_17, P0_17;
wire G0_18, P0_18;
wire G0_19, P0_19;
wire G0_20, P0_20;
wire G0_21, P0_21;
wire G0_22, P0_22;
wire G0_23, P0_23;
wire G0_24, P0_24;
wire G0_25, P0_25;
wire G0_26, P0_26;
wire G0_27, P0_27;
wire G0_28, P0_28;
wire G0_29, P0_29;
wire G0_30, P0_30;
wire G0_31, P0_31;
wire G0_32, P0_32;
wire G0_33, P0_33;
wire G0_34, P0_34;
wire G0_35, P0_35;
wire G0_36, P0_36;
wire G0_37, P0_37;
wire G0_38, P0_38;
wire G0_39, P0_39;
wire G0_40, P0_40;
wire G0_41, P0_41;
wire G0_42, P0_42;
wire G0_43, P0_43;
wire G0_44, P0_44;
wire G0_45, P0_45;
wire G0_46, P0_46;
wire G0_47, P0_47;
wire G0_48, P0_48;
wire G0_49, P0_49;
wire G0_50, P0_50;
wire G0_51, P0_51;
wire G0_52, P0_52;
wire G0_53, P0_53;
wire G0_54, P0_54;
wire G0_55, P0_55;
wire G0_56, P0_56;
wire G0_57, P0_57;
wire G0_58, P0_58;
wire G0_59, P0_59;
wire G0_60, P0_60;
wire G0_61, P0_61;
wire G0_62, P0_62;
wire G0_63, P0_63;
wire G1_0, P1_0;
wire G1_1, P1_1;
wire G1_2, P1_2;
wire G1_3, P1_3;
wire G1_4, P1_4;
wire G1_5, P1_5;
wire G1_6, P1_6;
wire G1_7, P1_7;
wire G1_8, P1_8;
wire G1_9, P1_9;
wire G1_10, P1_10;
wire G1_11, P1_11;
wire G1_12, P1_12;
wire G1_13, P1_13;
wire G1_14, P1_14;
wire G1_15, P1_15;
wire G1_16, P1_16;
wire G1_17, P1_17;
wire G1_18, P1_18;
wire G1_19, P1_19;
wire G1_20, P1_20;
wire G1_21, P1_21;
wire G1_22, P1_22;
wire G1_23, P1_23;
wire G1_24, P1_24;
wire G1_25, P1_25;
wire G1_26, P1_26;
wire G1_27, P1_27;
wire G1_28, P1_28;
wire G1_29, P1_29;
wire G1_30, P1_30;
wire G1_31, P1_31;
wire G1_32, P1_32;
wire G1_33, P1_33;
wire G1_34, P1_34;
wire G1_35, P1_35;
wire G1_36, P1_36;
wire G1_37, P1_37;
wire G1_38, P1_38;
wire G1_39, P1_39;
wire G1_40, P1_40;
wire G1_41, P1_41;
wire G1_42, P1_42;
wire G1_43, P1_43;
wire G1_44, P1_44;
wire G1_45, P1_45;
wire G1_46, P1_46;
wire G1_47, P1_47;
wire G1_48, P1_48;
wire G1_49, P1_49;
wire G1_50, P1_50;
wire G1_51, P1_51;
wire G1_52, P1_52;
wire G1_53, P1_53;
wire G1_54, P1_54;
wire G1_55, P1_55;
wire G1_56, P1_56;
wire G1_57, P1_57;
wire G1_58, P1_58;
wire G1_59, P1_59;
wire G1_60, P1_60;
wire G1_61, P1_61;
wire G1_62, P1_62;
wire G1_63, P1_63;
wire G2_0, P2_0;
wire G2_1, P2_1;
wire G2_2, P2_2;
wire G2_3, P2_3;
wire G2_4, P2_4;
wire G2_5, P2_5;
wire G2_6, P2_6;
wire G2_7, P2_7;
wire G2_8, P2_8;
wire G2_9, P2_9;
wire G2_10, P2_10;
wire G2_11, P2_11;
wire G2_12, P2_12;
wire G2_13, P2_13;
wire G2_14, P2_14;
wire G2_15, P2_15;
wire G2_16, P2_16;
wire G2_17, P2_17;
wire G2_18, P2_18;
wire G2_19, P2_19;
wire G2_20, P2_20;
wire G2_21, P2_21;
wire G2_22, P2_22;
wire G2_23, P2_23;
wire G2_24, P2_24;
wire G2_25, P2_25;
wire G2_26, P2_26;
wire G2_27, P2_27;
wire G2_28, P2_28;
wire G2_29, P2_29;
wire G2_30, P2_30;
wire G2_31, P2_31;
wire G2_32, P2_32;
wire G2_33, P2_33;
wire G2_34, P2_34;
wire G2_35, P2_35;
wire G2_36, P2_36;
wire G2_37, P2_37;
wire G2_38, P2_38;
wire G2_39, P2_39;
wire G2_40, P2_40;
wire G2_41, P2_41;
wire G2_42, P2_42;
wire G2_43, P2_43;
wire G2_44, P2_44;
wire G2_45, P2_45;
wire G2_46, P2_46;
wire G2_47, P2_47;
wire G2_48, P2_48;
wire G2_49, P2_49;
wire G2_50, P2_50;
wire G2_51, P2_51;
wire G2_52, P2_52;
wire G2_53, P2_53;
wire G2_54, P2_54;
wire G2_55, P2_55;
wire G2_56, P2_56;
wire G2_57, P2_57;
wire G2_58, P2_58;
wire G2_59, P2_59;
wire G2_60, P2_60;
wire G2_61, P2_61;
wire G2_62, P2_62;
wire G2_63, P2_63;
wire G3_0, P3_0;
wire G3_1, P3_1;
wire G3_2, P3_2;
wire G3_3, P3_3;
wire G3_4, P3_4;
wire G3_5, P3_5;
wire G3_6, P3_6;
wire G3_7, P3_7;
wire G3_8, P3_8;
wire G3_9, P3_9;
wire G3_10, P3_10;
wire G3_11, P3_11;
wire G3_12, P3_12;
wire G3_13, P3_13;
wire G3_14, P3_14;
wire G3_15, P3_15;
wire G3_16, P3_16;
wire G3_17, P3_17;
wire G3_18, P3_18;
wire G3_19, P3_19;
wire G3_20, P3_20;
wire G3_21, P3_21;
wire G3_22, P3_22;
wire G3_23, P3_23;
wire G3_24, P3_24;
wire G3_25, P3_25;
wire G3_26, P3_26;
wire G3_27, P3_27;
wire G3_28, P3_28;
wire G3_29, P3_29;
wire G3_30, P3_30;
wire G3_31, P3_31;
wire G3_32, P3_32;
wire G3_33, P3_33;
wire G3_34, P3_34;
wire G3_35, P3_35;
wire G3_36, P3_36;
wire G3_37, P3_37;
wire G3_38, P3_38;
wire G3_39, P3_39;
wire G3_40, P3_40;
wire G3_41, P3_41;
wire G3_42, P3_42;
wire G3_43, P3_43;
wire G3_44, P3_44;
wire G3_45, P3_45;
wire G3_46, P3_46;
wire G3_47, P3_47;
wire G3_48, P3_48;
wire G3_49, P3_49;
wire G3_50, P3_50;
wire G3_51, P3_51;
wire G3_52, P3_52;
wire G3_53, P3_53;
wire G3_54, P3_54;
wire G3_55, P3_55;
wire G3_56, P3_56;
wire G3_57, P3_57;
wire G3_58, P3_58;
wire G3_59, P3_59;
wire G3_60, P3_60;
wire G3_61, P3_61;
wire G3_62, P3_62;
wire G3_63, P3_63;
wire G4_0, P4_0;
wire G4_1, P4_1;
wire G4_2, P4_2;
wire G4_3, P4_3;
wire G4_4, P4_4;
wire G4_5, P4_5;
wire G4_6, P4_6;
wire G4_7, P4_7;
wire G4_8, P4_8;
wire G4_9, P4_9;
wire G4_10, P4_10;
wire G4_11, P4_11;
wire G4_12, P4_12;
wire G4_13, P4_13;
wire G4_14, P4_14;
wire G4_15, P4_15;
wire G4_16, P4_16;
wire G4_17, P4_17;
wire G4_18, P4_18;
wire G4_19, P4_19;
wire G4_20, P4_20;
wire G4_21, P4_21;
wire G4_22, P4_22;
wire G4_23, P4_23;
wire G4_24, P4_24;
wire G4_25, P4_25;
wire G4_26, P4_26;
wire G4_27, P4_27;
wire G4_28, P4_28;
wire G4_29, P4_29;
wire G4_30, P4_30;
wire G4_31, P4_31;
wire G4_32, P4_32;
wire G4_33, P4_33;
wire G4_34, P4_34;
wire G4_35, P4_35;
wire G4_36, P4_36;
wire G4_37, P4_37;
wire G4_38, P4_38;
wire G4_39, P4_39;
wire G4_40, P4_40;
wire G4_41, P4_41;
wire G4_42, P4_42;
wire G4_43, P4_43;
wire G4_44, P4_44;
wire G4_45, P4_45;
wire G4_46, P4_46;
wire G4_47, P4_47;
wire G4_48, P4_48;
wire G4_49, P4_49;
wire G4_50, P4_50;
wire G4_51, P4_51;
wire G4_52, P4_52;
wire G4_53, P4_53;
wire G4_54, P4_54;
wire G4_55, P4_55;
wire G4_56, P4_56;
wire G4_57, P4_57;
wire G4_58, P4_58;
wire G4_59, P4_59;
wire G4_60, P4_60;
wire G4_61, P4_61;
wire G4_62, P4_62;
wire G4_63, P4_63;
wire G5_0, P5_0;
wire G5_1, P5_1;
wire G5_2, P5_2;
wire G5_3, P5_3;
wire G5_4, P5_4;
wire G5_5, P5_5;
wire G5_6, P5_6;
wire G5_7, P5_7;
wire G5_8, P5_8;
wire G5_9, P5_9;
wire G5_10, P5_10;
wire G5_11, P5_11;
wire G5_12, P5_12;
wire G5_13, P5_13;
wire G5_14, P5_14;
wire G5_15, P5_15;
wire G5_16, P5_16;
wire G5_17, P5_17;
wire G5_18, P5_18;
wire G5_19, P5_19;
wire G5_20, P5_20;
wire G5_21, P5_21;
wire G5_22, P5_22;
wire G5_23, P5_23;
wire G5_24, P5_24;
wire G5_25, P5_25;
wire G5_26, P5_26;
wire G5_27, P5_27;
wire G5_28, P5_28;
wire G5_29, P5_29;
wire G5_30, P5_30;
wire G5_31, P5_31;
wire G5_32, P5_32;
wire G5_33, P5_33;
wire G5_34, P5_34;
wire G5_35, P5_35;
wire G5_36, P5_36;
wire G5_37, P5_37;
wire G5_38, P5_38;
wire G5_39, P5_39;
wire G5_40, P5_40;
wire G5_41, P5_41;
wire G5_42, P5_42;
wire G5_43, P5_43;
wire G5_44, P5_44;
wire G5_45, P5_45;
wire G5_46, P5_46;
wire G5_47, P5_47;
wire G5_48, P5_48;
wire G5_49, P5_49;
wire G5_50, P5_50;
wire G5_51, P5_51;
wire G5_52, P5_52;
wire G5_53, P5_53;
wire G5_54, P5_54;
wire G5_55, P5_55;
wire G5_56, P5_56;
wire G5_57, P5_57;
wire G5_58, P5_58;
wire G5_59, P5_59;
wire G5_60, P5_60;
wire G5_61, P5_61;
wire G5_62, P5_62;
wire G5_63, P5_63;

assign G0_0 = g[0];
assign P0_0 = p[0];
assign G0_1 = g[1];
assign P0_1 = p[1];
assign G0_2 = g[2];
assign P0_2 = p[2];
assign G0_3 = g[3];
assign P0_3 = p[3];
assign G0_4 = g[4];
assign P0_4 = p[4];
assign G0_5 = g[5];
assign P0_5 = p[5];
assign G0_6 = g[6];
assign P0_6 = p[6];
assign G0_7 = g[7];
assign P0_7 = p[7];
assign G0_8 = g[8];
assign P0_8 = p[8];
assign G0_9 = g[9];
assign P0_9 = p[9];
assign G0_10 = g[10];
assign P0_10 = p[10];
assign G0_11 = g[11];
assign P0_11 = p[11];
assign G0_12 = g[12];
assign P0_12 = p[12];
assign G0_13 = g[13];
assign P0_13 = p[13];
assign G0_14 = g[14];
assign P0_14 = p[14];
assign G0_15 = g[15];
assign P0_15 = p[15];
assign G0_16 = g[16];
assign P0_16 = p[16];
assign G0_17 = g[17];
assign P0_17 = p[17];
assign G0_18 = g[18];
assign P0_18 = p[18];
assign G0_19 = g[19];
assign P0_19 = p[19];
assign G0_20 = g[20];
assign P0_20 = p[20];
assign G0_21 = g[21];
assign P0_21 = p[21];
assign G0_22 = g[22];
assign P0_22 = p[22];
assign G0_23 = g[23];
assign P0_23 = p[23];
assign G0_24 = g[24];
assign P0_24 = p[24];
assign G0_25 = g[25];
assign P0_25 = p[25];
assign G0_26 = g[26];
assign P0_26 = p[26];
assign G0_27 = g[27];
assign P0_27 = p[27];
assign G0_28 = g[28];
assign P0_28 = p[28];
assign G0_29 = g[29];
assign P0_29 = p[29];
assign G0_30 = g[30];
assign P0_30 = p[30];
assign G0_31 = g[31];
assign P0_31 = p[31];
assign G0_32 = g[32];
assign P0_32 = p[32];
assign G0_33 = g[33];
assign P0_33 = p[33];
assign G0_34 = g[34];
assign P0_34 = p[34];
assign G0_35 = g[35];
assign P0_35 = p[35];
assign G0_36 = g[36];
assign P0_36 = p[36];
assign G0_37 = g[37];
assign P0_37 = p[37];
assign G0_38 = g[38];
assign P0_38 = p[38];
assign G0_39 = g[39];
assign P0_39 = p[39];
assign G0_40 = g[40];
assign P0_40 = p[40];
assign G0_41 = g[41];
assign P0_41 = p[41];
assign G0_42 = g[42];
assign P0_42 = p[42];
assign G0_43 = g[43];
assign P0_43 = p[43];
assign G0_44 = g[44];
assign P0_44 = p[44];
assign G0_45 = g[45];
assign P0_45 = p[45];
assign G0_46 = g[46];
assign P0_46 = p[46];
assign G0_47 = g[47];
assign P0_47 = p[47];
assign G0_48 = g[48];
assign P0_48 = p[48];
assign G0_49 = g[49];
assign P0_49 = p[49];
assign G0_50 = g[50];
assign P0_50 = p[50];
assign G0_51 = g[51];
assign P0_51 = p[51];
assign G0_52 = g[52];
assign P0_52 = p[52];
assign G0_53 = g[53];
assign P0_53 = p[53];
assign G0_54 = g[54];
assign P0_54 = p[54];
assign G0_55 = g[55];
assign P0_55 = p[55];
assign G0_56 = g[56];
assign P0_56 = p[56];
assign G0_57 = g[57];
assign P0_57 = p[57];
assign G0_58 = g[58];
assign P0_58 = p[58];
assign G0_59 = g[59];
assign P0_59 = p[59];
assign G0_60 = g[60];
assign P0_60 = p[60];
assign G0_61 = g[61];
assign P0_61 = p[61];
assign G0_62 = g[62];
assign P0_62 = p[62];
assign G0_63 = g[63];
assign P0_63 = p[63];

assign G1_0 = G0_0;
assign P1_0 = P0_0;
carry_operator s1_1 (G0_0, G0_1, P0_0, P0_1, G1_1, P1_1);
carry_operator s1_2 (G0_1, G0_2, P0_1, P0_2, G1_2, P1_2);
carry_operator s1_3 (G0_2, G0_3, P0_2, P0_3, G1_3, P1_3);
carry_operator s1_4 (G0_3, G0_4, P0_3, P0_4, G1_4, P1_4);
carry_operator s1_5 (G0_4, G0_5, P0_4, P0_5, G1_5, P1_5);
carry_operator s1_6 (G0_5, G0_6, P0_5, P0_6, G1_6, P1_6);
carry_operator s1_7 (G0_6, G0_7, P0_6, P0_7, G1_7, P1_7);
carry_operator s1_8 (G0_7, G0_8, P0_7, P0_8, G1_8, P1_8);
carry_operator s1_9 (G0_8, G0_9, P0_8, P0_9, G1_9, P1_9);
carry_operator s1_10 (G0_9, G0_10, P0_9, P0_10, G1_10, P1_10);
carry_operator s1_11 (G0_10, G0_11, P0_10, P0_11, G1_11, P1_11);
carry_operator s1_12 (G0_11, G0_12, P0_11, P0_12, G1_12, P1_12);
carry_operator s1_13 (G0_12, G0_13, P0_12, P0_13, G1_13, P1_13);
carry_operator s1_14 (G0_13, G0_14, P0_13, P0_14, G1_14, P1_14);
carry_operator s1_15 (G0_14, G0_15, P0_14, P0_15, G1_15, P1_15);
carry_operator s1_16 (G0_15, G0_16, P0_15, P0_16, G1_16, P1_16);
carry_operator s1_17 (G0_16, G0_17, P0_16, P0_17, G1_17, P1_17);
carry_operator s1_18 (G0_17, G0_18, P0_17, P0_18, G1_18, P1_18);
carry_operator s1_19 (G0_18, G0_19, P0_18, P0_19, G1_19, P1_19);
carry_operator s1_20 (G0_19, G0_20, P0_19, P0_20, G1_20, P1_20);
carry_operator s1_21 (G0_20, G0_21, P0_20, P0_21, G1_21, P1_21);
carry_operator s1_22 (G0_21, G0_22, P0_21, P0_22, G1_22, P1_22);
carry_operator s1_23 (G0_22, G0_23, P0_22, P0_23, G1_23, P1_23);
carry_operator s1_24 (G0_23, G0_24, P0_23, P0_24, G1_24, P1_24);
carry_operator s1_25 (G0_24, G0_25, P0_24, P0_25, G1_25, P1_25);
carry_operator s1_26 (G0_25, G0_26, P0_25, P0_26, G1_26, P1_26);
carry_operator s1_27 (G0_26, G0_27, P0_26, P0_27, G1_27, P1_27);
carry_operator s1_28 (G0_27, G0_28, P0_27, P0_28, G1_28, P1_28);
carry_operator s1_29 (G0_28, G0_29, P0_28, P0_29, G1_29, P1_29);
carry_operator s1_30 (G0_29, G0_30, P0_29, P0_30, G1_30, P1_30);
carry_operator s1_31 (G0_30, G0_31, P0_30, P0_31, G1_31, P1_31);
carry_operator s1_32 (G0_31, G0_32, P0_31, P0_32, G1_32, P1_32);
carry_operator s1_33 (G0_32, G0_33, P0_32, P0_33, G1_33, P1_33);
carry_operator s1_34 (G0_33, G0_34, P0_33, P0_34, G1_34, P1_34);
carry_operator s1_35 (G0_34, G0_35, P0_34, P0_35, G1_35, P1_35);
carry_operator s1_36 (G0_35, G0_36, P0_35, P0_36, G1_36, P1_36);
carry_operator s1_37 (G0_36, G0_37, P0_36, P0_37, G1_37, P1_37);
carry_operator s1_38 (G0_37, G0_38, P0_37, P0_38, G1_38, P1_38);
carry_operator s1_39 (G0_38, G0_39, P0_38, P0_39, G1_39, P1_39);
carry_operator s1_40 (G0_39, G0_40, P0_39, P0_40, G1_40, P1_40);
carry_operator s1_41 (G0_40, G0_41, P0_40, P0_41, G1_41, P1_41);
carry_operator s1_42 (G0_41, G0_42, P0_41, P0_42, G1_42, P1_42);
carry_operator s1_43 (G0_42, G0_43, P0_42, P0_43, G1_43, P1_43);
carry_operator s1_44 (G0_43, G0_44, P0_43, P0_44, G1_44, P1_44);
carry_operator s1_45 (G0_44, G0_45, P0_44, P0_45, G1_45, P1_45);
carry_operator s1_46 (G0_45, G0_46, P0_45, P0_46, G1_46, P1_46);
carry_operator s1_47 (G0_46, G0_47, P0_46, P0_47, G1_47, P1_47);
carry_operator s1_48 (G0_47, G0_48, P0_47, P0_48, G1_48, P1_48);
carry_operator s1_49 (G0_48, G0_49, P0_48, P0_49, G1_49, P1_49);
carry_operator s1_50 (G0_49, G0_50, P0_49, P0_50, G1_50, P1_50);
carry_operator s1_51 (G0_50, G0_51, P0_50, P0_51, G1_51, P1_51);
carry_operator s1_52 (G0_51, G0_52, P0_51, P0_52, G1_52, P1_52);
carry_operator s1_53 (G0_52, G0_53, P0_52, P0_53, G1_53, P1_53);
carry_operator s1_54 (G0_53, G0_54, P0_53, P0_54, G1_54, P1_54);
carry_operator s1_55 (G0_54, G0_55, P0_54, P0_55, G1_55, P1_55);
carry_operator s1_56 (G0_55, G0_56, P0_55, P0_56, G1_56, P1_56);
carry_operator s1_57 (G0_56, G0_57, P0_56, P0_57, G1_57, P1_57);
carry_operator s1_58 (G0_57, G0_58, P0_57, P0_58, G1_58, P1_58);
carry_operator s1_59 (G0_58, G0_59, P0_58, P0_59, G1_59, P1_59);
carry_operator s1_60 (G0_59, G0_60, P0_59, P0_60, G1_60, P1_60);
carry_operator s1_61 (G0_60, G0_61, P0_60, P0_61, G1_61, P1_61);
carry_operator s1_62 (G0_61, G0_62, P0_61, P0_62, G1_62, P1_62);
carry_operator s1_63 (G0_62, G0_63, P0_62, P0_63, G1_63, P1_63);

assign G2_0 = G1_0;
assign P2_0 = P1_0;
assign G2_1 = G1_1;
assign P2_1 = P1_1;
carry_operator s2_2 (G1_0, G1_2, P1_0, P1_2, G2_2, P2_2);
carry_operator s2_3 (G1_1, G1_3, P1_1, P1_3, G2_3, P2_3);
carry_operator s2_4 (G1_2, G1_4, P1_2, P1_4, G2_4, P2_4);
carry_operator s2_5 (G1_3, G1_5, P1_3, P1_5, G2_5, P2_5);
carry_operator s2_6 (G1_4, G1_6, P1_4, P1_6, G2_6, P2_6);
carry_operator s2_7 (G1_5, G1_7, P1_5, P1_7, G2_7, P2_7);
carry_operator s2_8 (G1_6, G1_8, P1_6, P1_8, G2_8, P2_8);
carry_operator s2_9 (G1_7, G1_9, P1_7, P1_9, G2_9, P2_9);
carry_operator s2_10 (G1_8, G1_10, P1_8, P1_10, G2_10, P2_10);
carry_operator s2_11 (G1_9, G1_11, P1_9, P1_11, G2_11, P2_11);
carry_operator s2_12 (G1_10, G1_12, P1_10, P1_12, G2_12, P2_12);
carry_operator s2_13 (G1_11, G1_13, P1_11, P1_13, G2_13, P2_13);
carry_operator s2_14 (G1_12, G1_14, P1_12, P1_14, G2_14, P2_14);
carry_operator s2_15 (G1_13, G1_15, P1_13, P1_15, G2_15, P2_15);
carry_operator s2_16 (G1_14, G1_16, P1_14, P1_16, G2_16, P2_16);
carry_operator s2_17 (G1_15, G1_17, P1_15, P1_17, G2_17, P2_17);
carry_operator s2_18 (G1_16, G1_18, P1_16, P1_18, G2_18, P2_18);
carry_operator s2_19 (G1_17, G1_19, P1_17, P1_19, G2_19, P2_19);
carry_operator s2_20 (G1_18, G1_20, P1_18, P1_20, G2_20, P2_20);
carry_operator s2_21 (G1_19, G1_21, P1_19, P1_21, G2_21, P2_21);
carry_operator s2_22 (G1_20, G1_22, P1_20, P1_22, G2_22, P2_22);
carry_operator s2_23 (G1_21, G1_23, P1_21, P1_23, G2_23, P2_23);
carry_operator s2_24 (G1_22, G1_24, P1_22, P1_24, G2_24, P2_24);
carry_operator s2_25 (G1_23, G1_25, P1_23, P1_25, G2_25, P2_25);
carry_operator s2_26 (G1_24, G1_26, P1_24, P1_26, G2_26, P2_26);
carry_operator s2_27 (G1_25, G1_27, P1_25, P1_27, G2_27, P2_27);
carry_operator s2_28 (G1_26, G1_28, P1_26, P1_28, G2_28, P2_28);
carry_operator s2_29 (G1_27, G1_29, P1_27, P1_29, G2_29, P2_29);
carry_operator s2_30 (G1_28, G1_30, P1_28, P1_30, G2_30, P2_30);
carry_operator s2_31 (G1_29, G1_31, P1_29, P1_31, G2_31, P2_31);
carry_operator s2_32 (G1_30, G1_32, P1_30, P1_32, G2_32, P2_32);
carry_operator s2_33 (G1_31, G1_33, P1_31, P1_33, G2_33, P2_33);
carry_operator s2_34 (G1_32, G1_34, P1_32, P1_34, G2_34, P2_34);
carry_operator s2_35 (G1_33, G1_35, P1_33, P1_35, G2_35, P2_35);
carry_operator s2_36 (G1_34, G1_36, P1_34, P1_36, G2_36, P2_36);
carry_operator s2_37 (G1_35, G1_37, P1_35, P1_37, G2_37, P2_37);
carry_operator s2_38 (G1_36, G1_38, P1_36, P1_38, G2_38, P2_38);
carry_operator s2_39 (G1_37, G1_39, P1_37, P1_39, G2_39, P2_39);
carry_operator s2_40 (G1_38, G1_40, P1_38, P1_40, G2_40, P2_40);
carry_operator s2_41 (G1_39, G1_41, P1_39, P1_41, G2_41, P2_41);
carry_operator s2_42 (G1_40, G1_42, P1_40, P1_42, G2_42, P2_42);
carry_operator s2_43 (G1_41, G1_43, P1_41, P1_43, G2_43, P2_43);
carry_operator s2_44 (G1_42, G1_44, P1_42, P1_44, G2_44, P2_44);
carry_operator s2_45 (G1_43, G1_45, P1_43, P1_45, G2_45, P2_45);
carry_operator s2_46 (G1_44, G1_46, P1_44, P1_46, G2_46, P2_46);
carry_operator s2_47 (G1_45, G1_47, P1_45, P1_47, G2_47, P2_47);
carry_operator s2_48 (G1_46, G1_48, P1_46, P1_48, G2_48, P2_48);
carry_operator s2_49 (G1_47, G1_49, P1_47, P1_49, G2_49, P2_49);
carry_operator s2_50 (G1_48, G1_50, P1_48, P1_50, G2_50, P2_50);
carry_operator s2_51 (G1_49, G1_51, P1_49, P1_51, G2_51, P2_51);
carry_operator s2_52 (G1_50, G1_52, P1_50, P1_52, G2_52, P2_52);
carry_operator s2_53 (G1_51, G1_53, P1_51, P1_53, G2_53, P2_53);
carry_operator s2_54 (G1_52, G1_54, P1_52, P1_54, G2_54, P2_54);
carry_operator s2_55 (G1_53, G1_55, P1_53, P1_55, G2_55, P2_55);
carry_operator s2_56 (G1_54, G1_56, P1_54, P1_56, G2_56, P2_56);
carry_operator s2_57 (G1_55, G1_57, P1_55, P1_57, G2_57, P2_57);
carry_operator s2_58 (G1_56, G1_58, P1_56, P1_58, G2_58, P2_58);
carry_operator s2_59 (G1_57, G1_59, P1_57, P1_59, G2_59, P2_59);
carry_operator s2_60 (G1_58, G1_60, P1_58, P1_60, G2_60, P2_60);
carry_operator s2_61 (G1_59, G1_61, P1_59, P1_61, G2_61, P2_61);
carry_operator s2_62 (G1_60, G1_62, P1_60, P1_62, G2_62, P2_62);
carry_operator s2_63 (G1_61, G1_63, P1_61, P1_63, G2_63, P2_63);

assign G3_0 = G2_0;
assign P3_0 = P2_0;
assign G3_1 = G2_1;
assign P3_1 = P2_1;
assign G3_2 = G2_2;
assign P3_2 = P2_2;
assign G3_3 = G2_3;
assign P3_3 = P2_3;
carry_operator s3_4 (G2_0, G2_4, P2_0, P2_4, G3_4, P3_4);
carry_operator s3_5 (G2_1, G2_5, P2_1, P2_5, G3_5, P3_5);
carry_operator s3_6 (G2_2, G2_6, P2_2, P2_6, G3_6, P3_6);
carry_operator s3_7 (G2_3, G2_7, P2_3, P2_7, G3_7, P3_7);
carry_operator s3_8 (G2_4, G2_8, P2_4, P2_8, G3_8, P3_8);
carry_operator s3_9 (G2_5, G2_9, P2_5, P2_9, G3_9, P3_9);
carry_operator s3_10 (G2_6, G2_10, P2_6, P2_10, G3_10, P3_10);
carry_operator s3_11 (G2_7, G2_11, P2_7, P2_11, G3_11, P3_11);
carry_operator s3_12 (G2_8, G2_12, P2_8, P2_12, G3_12, P3_12);
carry_operator s3_13 (G2_9, G2_13, P2_9, P2_13, G3_13, P3_13);
carry_operator s3_14 (G2_10, G2_14, P2_10, P2_14, G3_14, P3_14);
carry_operator s3_15 (G2_11, G2_15, P2_11, P2_15, G3_15, P3_15);
carry_operator s3_16 (G2_12, G2_16, P2_12, P2_16, G3_16, P3_16);
carry_operator s3_17 (G2_13, G2_17, P2_13, P2_17, G3_17, P3_17);
carry_operator s3_18 (G2_14, G2_18, P2_14, P2_18, G3_18, P3_18);
carry_operator s3_19 (G2_15, G2_19, P2_15, P2_19, G3_19, P3_19);
carry_operator s3_20 (G2_16, G2_20, P2_16, P2_20, G3_20, P3_20);
carry_operator s3_21 (G2_17, G2_21, P2_17, P2_21, G3_21, P3_21);
carry_operator s3_22 (G2_18, G2_22, P2_18, P2_22, G3_22, P3_22);
carry_operator s3_23 (G2_19, G2_23, P2_19, P2_23, G3_23, P3_23);
carry_operator s3_24 (G2_20, G2_24, P2_20, P2_24, G3_24, P3_24);
carry_operator s3_25 (G2_21, G2_25, P2_21, P2_25, G3_25, P3_25);
carry_operator s3_26 (G2_22, G2_26, P2_22, P2_26, G3_26, P3_26);
carry_operator s3_27 (G2_23, G2_27, P2_23, P2_27, G3_27, P3_27);
carry_operator s3_28 (G2_24, G2_28, P2_24, P2_28, G3_28, P3_28);
carry_operator s3_29 (G2_25, G2_29, P2_25, P2_29, G3_29, P3_29);
carry_operator s3_30 (G2_26, G2_30, P2_26, P2_30, G3_30, P3_30);
carry_operator s3_31 (G2_27, G2_31, P2_27, P2_31, G3_31, P3_31);
carry_operator s3_32 (G2_28, G2_32, P2_28, P2_32, G3_32, P3_32);
carry_operator s3_33 (G2_29, G2_33, P2_29, P2_33, G3_33, P3_33);
carry_operator s3_34 (G2_30, G2_34, P2_30, P2_34, G3_34, P3_34);
carry_operator s3_35 (G2_31, G2_35, P2_31, P2_35, G3_35, P3_35);
carry_operator s3_36 (G2_32, G2_36, P2_32, P2_36, G3_36, P3_36);
carry_operator s3_37 (G2_33, G2_37, P2_33, P2_37, G3_37, P3_37);
carry_operator s3_38 (G2_34, G2_38, P2_34, P2_38, G3_38, P3_38);
carry_operator s3_39 (G2_35, G2_39, P2_35, P2_39, G3_39, P3_39);
carry_operator s3_40 (G2_36, G2_40, P2_36, P2_40, G3_40, P3_40);
carry_operator s3_41 (G2_37, G2_41, P2_37, P2_41, G3_41, P3_41);
carry_operator s3_42 (G2_38, G2_42, P2_38, P2_42, G3_42, P3_42);
carry_operator s3_43 (G2_39, G2_43, P2_39, P2_43, G3_43, P3_43);
carry_operator s3_44 (G2_40, G2_44, P2_40, P2_44, G3_44, P3_44);
carry_operator s3_45 (G2_41, G2_45, P2_41, P2_45, G3_45, P3_45);
carry_operator s3_46 (G2_42, G2_46, P2_42, P2_46, G3_46, P3_46);
carry_operator s3_47 (G2_43, G2_47, P2_43, P2_47, G3_47, P3_47);
carry_operator s3_48 (G2_44, G2_48, P2_44, P2_48, G3_48, P3_48);
carry_operator s3_49 (G2_45, G2_49, P2_45, P2_49, G3_49, P3_49);
carry_operator s3_50 (G2_46, G2_50, P2_46, P2_50, G3_50, P3_50);
carry_operator s3_51 (G2_47, G2_51, P2_47, P2_51, G3_51, P3_51);
carry_operator s3_52 (G2_48, G2_52, P2_48, P2_52, G3_52, P3_52);
carry_operator s3_53 (G2_49, G2_53, P2_49, P2_53, G3_53, P3_53);
carry_operator s3_54 (G2_50, G2_54, P2_50, P2_54, G3_54, P3_54);
carry_operator s3_55 (G2_51, G2_55, P2_51, P2_55, G3_55, P3_55);
carry_operator s3_56 (G2_52, G2_56, P2_52, P2_56, G3_56, P3_56);
carry_operator s3_57 (G2_53, G2_57, P2_53, P2_57, G3_57, P3_57);
carry_operator s3_58 (G2_54, G2_58, P2_54, P2_58, G3_58, P3_58);
carry_operator s3_59 (G2_55, G2_59, P2_55, P2_59, G3_59, P3_59);
carry_operator s3_60 (G2_56, G2_60, P2_56, P2_60, G3_60, P3_60);
carry_operator s3_61 (G2_57, G2_61, P2_57, P2_61, G3_61, P3_61);
carry_operator s3_62 (G2_58, G2_62, P2_58, P2_62, G3_62, P3_62);
carry_operator s3_63 (G2_59, G2_63, P2_59, P2_63, G3_63, P3_63);

assign G4_0 = G3_0;
assign P4_0 = P3_0;
assign G4_1 = G3_1;
assign P4_1 = P3_1;
assign G4_2 = G3_2;
assign P4_2 = P3_2;
assign G4_3 = G3_3;
assign P4_3 = P3_3;
assign G4_4 = G3_4;
assign P4_4 = P3_4;
assign G4_5 = G3_5;
assign P4_5 = P3_5;
assign G4_6 = G3_6;
assign P4_6 = P3_6;
assign G4_7 = G3_7;
assign P4_7 = P3_7;
carry_operator s4_8 (G3_0, G3_8, P3_0, P3_8, G4_8, P4_8);
carry_operator s4_9 (G3_1, G3_9, P3_1, P3_9, G4_9, P4_9);
carry_operator s4_10 (G3_2, G3_10, P3_2, P3_10, G4_10, P4_10);
carry_operator s4_11 (G3_3, G3_11, P3_3, P3_11, G4_11, P4_11);
carry_operator s4_12 (G3_4, G3_12, P3_4, P3_12, G4_12, P4_12);
carry_operator s4_13 (G3_5, G3_13, P3_5, P3_13, G4_13, P4_13);
carry_operator s4_14 (G3_6, G3_14, P3_6, P3_14, G4_14, P4_14);
carry_operator s4_15 (G3_7, G3_15, P3_7, P3_15, G4_15, P4_15);
carry_operator s4_16 (G3_8, G3_16, P3_8, P3_16, G4_16, P4_16);
carry_operator s4_17 (G3_9, G3_17, P3_9, P3_17, G4_17, P4_17);
carry_operator s4_18 (G3_10, G3_18, P3_10, P3_18, G4_18, P4_18);
carry_operator s4_19 (G3_11, G3_19, P3_11, P3_19, G4_19, P4_19);
carry_operator s4_20 (G3_12, G3_20, P3_12, P3_20, G4_20, P4_20);
carry_operator s4_21 (G3_13, G3_21, P3_13, P3_21, G4_21, P4_21);
carry_operator s4_22 (G3_14, G3_22, P3_14, P3_22, G4_22, P4_22);
carry_operator s4_23 (G3_15, G3_23, P3_15, P3_23, G4_23, P4_23);
carry_operator s4_24 (G3_16, G3_24, P3_16, P3_24, G4_24, P4_24);
carry_operator s4_25 (G3_17, G3_25, P3_17, P3_25, G4_25, P4_25);
carry_operator s4_26 (G3_18, G3_26, P3_18, P3_26, G4_26, P4_26);
carry_operator s4_27 (G3_19, G3_27, P3_19, P3_27, G4_27, P4_27);
carry_operator s4_28 (G3_20, G3_28, P3_20, P3_28, G4_28, P4_28);
carry_operator s4_29 (G3_21, G3_29, P3_21, P3_29, G4_29, P4_29);
carry_operator s4_30 (G3_22, G3_30, P3_22, P3_30, G4_30, P4_30);
carry_operator s4_31 (G3_23, G3_31, P3_23, P3_31, G4_31, P4_31);
carry_operator s4_32 (G3_24, G3_32, P3_24, P3_32, G4_32, P4_32);
carry_operator s4_33 (G3_25, G3_33, P3_25, P3_33, G4_33, P4_33);
carry_operator s4_34 (G3_26, G3_34, P3_26, P3_34, G4_34, P4_34);
carry_operator s4_35 (G3_27, G3_35, P3_27, P3_35, G4_35, P4_35);
carry_operator s4_36 (G3_28, G3_36, P3_28, P3_36, G4_36, P4_36);
carry_operator s4_37 (G3_29, G3_37, P3_29, P3_37, G4_37, P4_37);
carry_operator s4_38 (G3_30, G3_38, P3_30, P3_38, G4_38, P4_38);
carry_operator s4_39 (G3_31, G3_39, P3_31, P3_39, G4_39, P4_39);
carry_operator s4_40 (G3_32, G3_40, P3_32, P3_40, G4_40, P4_40);
carry_operator s4_41 (G3_33, G3_41, P3_33, P3_41, G4_41, P4_41);
carry_operator s4_42 (G3_34, G3_42, P3_34, P3_42, G4_42, P4_42);
carry_operator s4_43 (G3_35, G3_43, P3_35, P3_43, G4_43, P4_43);
carry_operator s4_44 (G3_36, G3_44, P3_36, P3_44, G4_44, P4_44);
carry_operator s4_45 (G3_37, G3_45, P3_37, P3_45, G4_45, P4_45);
carry_operator s4_46 (G3_38, G3_46, P3_38, P3_46, G4_46, P4_46);
carry_operator s4_47 (G3_39, G3_47, P3_39, P3_47, G4_47, P4_47);
carry_operator s4_48 (G3_40, G3_48, P3_40, P3_48, G4_48, P4_48);
carry_operator s4_49 (G3_41, G3_49, P3_41, P3_49, G4_49, P4_49);
carry_operator s4_50 (G3_42, G3_50, P3_42, P3_50, G4_50, P4_50);
carry_operator s4_51 (G3_43, G3_51, P3_43, P3_51, G4_51, P4_51);
carry_operator s4_52 (G3_44, G3_52, P3_44, P3_52, G4_52, P4_52);
carry_operator s4_53 (G3_45, G3_53, P3_45, P3_53, G4_53, P4_53);
carry_operator s4_54 (G3_46, G3_54, P3_46, P3_54, G4_54, P4_54);
carry_operator s4_55 (G3_47, G3_55, P3_47, P3_55, G4_55, P4_55);
carry_operator s4_56 (G3_48, G3_56, P3_48, P3_56, G4_56, P4_56);
carry_operator s4_57 (G3_49, G3_57, P3_49, P3_57, G4_57, P4_57);
carry_operator s4_58 (G3_50, G3_58, P3_50, P3_58, G4_58, P4_58);
carry_operator s4_59 (G3_51, G3_59, P3_51, P3_59, G4_59, P4_59);
carry_operator s4_60 (G3_52, G3_60, P3_52, P3_60, G4_60, P4_60);
carry_operator s4_61 (G3_53, G3_61, P3_53, P3_61, G4_61, P4_61);
carry_operator s4_62 (G3_54, G3_62, P3_54, P3_62, G4_62, P4_62);
carry_operator s4_63 (G3_55, G3_63, P3_55, P3_63, G4_63, P4_63);

assign G5_0 = G4_0;
assign P5_0 = P4_0;
assign G5_1 = G4_1;
assign P5_1 = P4_1;
assign G5_2 = G4_2;
assign P5_2 = P4_2;
assign G5_3 = G4_3;
assign P5_3 = P4_3;
assign G5_4 = G4_4;
assign P5_4 = P4_4;
assign G5_5 = G4_5;
assign P5_5 = P4_5;
assign G5_6 = G4_6;
assign P5_6 = P4_6;
assign G5_7 = G4_7;
assign P5_7 = P4_7;
assign G5_8 = G4_8;
assign P5_8 = P4_8;
assign G5_9 = G4_9;
assign P5_9 = P4_9;
assign G5_10 = G4_10;
assign P5_10 = P4_10;
assign G5_11 = G4_11;
assign P5_11 = P4_11;
assign G5_12 = G4_12;
assign P5_12 = P4_12;
assign G5_13 = G4_13;
assign P5_13 = P4_13;
assign G5_14 = G4_14;
assign P5_14 = P4_14;
assign G5_15 = G4_15;
assign P5_15 = P4_15;
carry_operator s5_16 (G4_0, G4_16, P4_0, P4_16, G5_16, P5_16);
carry_operator s5_17 (G4_1, G4_17, P4_1, P4_17, G5_17, P5_17);
carry_operator s5_18 (G4_2, G4_18, P4_2, P4_18, G5_18, P5_18);
carry_operator s5_19 (G4_3, G4_19, P4_3, P4_19, G5_19, P5_19);
carry_operator s5_20 (G4_4, G4_20, P4_4, P4_20, G5_20, P5_20);
carry_operator s5_21 (G4_5, G4_21, P4_5, P4_21, G5_21, P5_21);
carry_operator s5_22 (G4_6, G4_22, P4_6, P4_22, G5_22, P5_22);
carry_operator s5_23 (G4_7, G4_23, P4_7, P4_23, G5_23, P5_23);
carry_operator s5_24 (G4_8, G4_24, P4_8, P4_24, G5_24, P5_24);
carry_operator s5_25 (G4_9, G4_25, P4_9, P4_25, G5_25, P5_25);
carry_operator s5_26 (G4_10, G4_26, P4_10, P4_26, G5_26, P5_26);
carry_operator s5_27 (G4_11, G4_27, P4_11, P4_27, G5_27, P5_27);
carry_operator s5_28 (G4_12, G4_28, P4_12, P4_28, G5_28, P5_28);
carry_operator s5_29 (G4_13, G4_29, P4_13, P4_29, G5_29, P5_29);
carry_operator s5_30 (G4_14, G4_30, P4_14, P4_30, G5_30, P5_30);
carry_operator s5_31 (G4_15, G4_31, P4_15, P4_31, G5_31, P5_31);
carry_operator s5_32 (G4_16, G4_32, P4_16, P4_32, G5_32, P5_32);
carry_operator s5_33 (G4_17, G4_33, P4_17, P4_33, G5_33, P5_33);
carry_operator s5_34 (G4_18, G4_34, P4_18, P4_34, G5_34, P5_34);
carry_operator s5_35 (G4_19, G4_35, P4_19, P4_35, G5_35, P5_35);
carry_operator s5_36 (G4_20, G4_36, P4_20, P4_36, G5_36, P5_36);
carry_operator s5_37 (G4_21, G4_37, P4_21, P4_37, G5_37, P5_37);
carry_operator s5_38 (G4_22, G4_38, P4_22, P4_38, G5_38, P5_38);
carry_operator s5_39 (G4_23, G4_39, P4_23, P4_39, G5_39, P5_39);
carry_operator s5_40 (G4_24, G4_40, P4_24, P4_40, G5_40, P5_40);
carry_operator s5_41 (G4_25, G4_41, P4_25, P4_41, G5_41, P5_41);
carry_operator s5_42 (G4_26, G4_42, P4_26, P4_42, G5_42, P5_42);
carry_operator s5_43 (G4_27, G4_43, P4_27, P4_43, G5_43, P5_43);
carry_operator s5_44 (G4_28, G4_44, P4_28, P4_44, G5_44, P5_44);
carry_operator s5_45 (G4_29, G4_45, P4_29, P4_45, G5_45, P5_45);
carry_operator s5_46 (G4_30, G4_46, P4_30, P4_46, G5_46, P5_46);
carry_operator s5_47 (G4_31, G4_47, P4_31, P4_47, G5_47, P5_47);
carry_operator s5_48 (G4_32, G4_48, P4_32, P4_48, G5_48, P5_48);
carry_operator s5_49 (G4_33, G4_49, P4_33, P4_49, G5_49, P5_49);
carry_operator s5_50 (G4_34, G4_50, P4_34, P4_50, G5_50, P5_50);
carry_operator s5_51 (G4_35, G4_51, P4_35, P4_51, G5_51, P5_51);
carry_operator s5_52 (G4_36, G4_52, P4_36, P4_52, G5_52, P5_52);
carry_operator s5_53 (G4_37, G4_53, P4_37, P4_53, G5_53, P5_53);
carry_operator s5_54 (G4_38, G4_54, P4_38, P4_54, G5_54, P5_54);
carry_operator s5_55 (G4_39, G4_55, P4_39, P4_55, G5_55, P5_55);
carry_operator s5_56 (G4_40, G4_56, P4_40, P4_56, G5_56, P5_56);
carry_operator s5_57 (G4_41, G4_57, P4_41, P4_57, G5_57, P5_57);
carry_operator s5_58 (G4_42, G4_58, P4_42, P4_58, G5_58, P5_58);
carry_operator s5_59 (G4_43, G4_59, P4_43, P4_59, G5_59, P5_59);
carry_operator s5_60 (G4_44, G4_60, P4_44, P4_60, G5_60, P5_60);
carry_operator s5_61 (G4_45, G4_61, P4_45, P4_61, G5_61, P5_61);
carry_operator s5_62 (G4_46, G4_62, P4_46, P4_62, G5_62, P5_62);
carry_operator s5_63 (G4_47, G4_63, P4_47, P4_63, G5_63, P5_63);

assign C[1] = G5_0 | (P5_0 & C[0]);
assign C[2] = G5_1 | (P5_1 & C[1]);
assign C[3] = G5_2 | (P5_2 & C[2]);
assign C[4] = G5_3 | (P5_3 & C[3]);
assign C[5] = G5_4 | (P5_4 & C[4]);
assign C[6] = G5_5 | (P5_5 & C[5]);
assign C[7] = G5_6 | (P5_6 & C[6]);
assign C[8] = G5_7 | (P5_7 & C[7]);
assign C[9] = G5_8 | (P5_8 & C[8]);
assign C[10] = G5_9 | (P5_9 & C[9]);
assign C[11] = G5_10 | (P5_10 & C[10]);
assign C[12] = G5_11 | (P5_11 & C[11]);
assign C[13] = G5_12 | (P5_12 & C[12]);
assign C[14] = G5_13 | (P5_13 & C[13]);
assign C[15] = G5_14 | (P5_14 & C[14]);
assign C[16] = G5_15 | (P5_15 & C[15]);
assign C[17] = G5_16 | (P5_16 & C[16]);
assign C[18] = G5_17 | (P5_17 & C[17]);
assign C[19] = G5_18 | (P5_18 & C[18]);
assign C[20] = G5_19 | (P5_19 & C[19]);
assign C[21] = G5_20 | (P5_20 & C[20]);
assign C[22] = G5_21 | (P5_21 & C[21]);
assign C[23] = G5_22 | (P5_22 & C[22]);
assign C[24] = G5_23 | (P5_23 & C[23]);
assign C[25] = G5_24 | (P5_24 & C[24]);
assign C[26] = G5_25 | (P5_25 & C[25]);
assign C[27] = G5_26 | (P5_26 & C[26]);
assign C[28] = G5_27 | (P5_27 & C[27]);
assign C[29] = G5_28 | (P5_28 & C[28]);
assign C[30] = G5_29 | (P5_29 & C[29]);
assign C[31] = G5_30 | (P5_30 & C[30]);
assign C[32] = G5_31 | (P5_31 & C[31]);
assign C[33] = G5_32 | (P5_32 & C[32]);
assign C[34] = G5_33 | (P5_33 & C[33]);
assign C[35] = G5_34 | (P5_34 & C[34]);
assign C[36] = G5_35 | (P5_35 & C[35]);
assign C[37] = G5_36 | (P5_36 & C[36]);
assign C[38] = G5_37 | (P5_37 & C[37]);
assign C[39] = G5_38 | (P5_38 & C[38]);
assign C[40] = G5_39 | (P5_39 & C[39]);
assign C[41] = G5_40 | (P5_40 & C[40]);
assign C[42] = G5_41 | (P5_41 & C[41]);
assign C[43] = G5_42 | (P5_42 & C[42]);
assign C[44] = G5_43 | (P5_43 & C[43]);
assign C[45] = G5_44 | (P5_44 & C[44]);
assign C[46] = G5_45 | (P5_45 & C[45]);
assign C[47] = G5_46 | (P5_46 & C[46]);
assign C[48] = G5_47 | (P5_47 & C[47]);
assign C[49] = G5_48 | (P5_48 & C[48]);
assign C[50] = G5_49 | (P5_49 & C[49]);
assign C[51] = G5_50 | (P5_50 & C[50]);
assign C[52] = G5_51 | (P5_51 & C[51]);
assign C[53] = G5_52 | (P5_52 & C[52]);
assign C[54] = G5_53 | (P5_53 & C[53]);
assign C[55] = G5_54 | (P5_54 & C[54]);
assign C[56] = G5_55 | (P5_55 & C[55]);
assign C[57] = G5_56 | (P5_56 & C[56]);
assign C[58] = G5_57 | (P5_57 & C[57]);
assign C[59] = G5_58 | (P5_58 & C[58]);
assign C[60] = G5_59 | (P5_59 & C[59]);
assign C[61] = G5_60 | (P5_60 & C[60]);
assign C[62] = G5_61 | (P5_61 & C[61]);
assign C[63] = G5_62 | (P5_62 & C[62]);
assign C[64] = G5_63 | (P5_63 & C[63]);
assign cout = C[64];
genvar i;
 generate
        for (i = 0; i < 64; i = i + 1) begin
            assign sum[i] = p[i] ^ C[i];
        end
    endgenerate

endmodule